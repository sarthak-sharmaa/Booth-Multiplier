module xor2 (
            input wire x, y, 
            output wire z
            );
  assign z = x ^ y;
endmodule
